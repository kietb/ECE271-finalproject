module sinWave (input logic s_clk,
		output logic [7:0] wave);

logic [9:0] count = 0;

always_ff @ (posedge s_clk) begin
  if (count >= 500)
    count <= 0;
    else 
      count <= count + 1;
end

always @(s_clk) begin
  case(count)

	0: wave <=127;
	1: wave <=129;
	2: wave <=130;
	3: wave <=132;
	4: wave <=133;
	5: wave <=135;	
	6: wave <=136;
	7: wave <=138;
	8: wave <=139;
	9: wave <=141;
	10: wave <=142;
	11: wave <=144;
	12: wave <=145;
	13: wave <=147;
	14: wave <=148;
	15: wave <=150;
	16: wave <=151;
	17: wave <=153;
	18: wave <=154;
	19: wave <=156;
	20: wave <=157;
	21: wave <=159;
	22: wave <=160;
	23: wave <=162;
	24: wave <=163;
	25: wave <=165;
	26: wave <=166;
	27: wave <=167;
	28: wave <=169;
	29: wave <=170;
	30: wave <=172;
31: wave <=173;
32: wave <=175;
33: wave <=176;
34: wave <=177;
35: wave <=179;
36: wave <=180;
37: wave <=182;
38: wave <=183;
39: wave <=184;
40: wave <=186;
41: wave <=187;
42: wave <=188;
43: wave <=190;
44: wave <=191;
45: wave <=192;
46: wave <=194;
47: wave <=195;
48: wave <=196;
49: wave <=198;
50: wave <=199;
51: wave <=200;
52: wave <=201;
53: wave <=203;
54: wave <=204;
55: wave <=205;
56: wave <=206;
57: wave <=207;
58: wave <=209;
59: wave <=210;
60: wave <=211;
61: wave <=212;
62: wave <=213;
63: wave <=214;
64: wave <=215;
65: wave <=216;
66: wave <=218;
67: wave <=219;
68: wave <=220;
69: wave <=221;
70: wave <=222;
71: wave <=223;
72: wave <=224;
73: wave <=225;
74: wave <=226;
75: wave <=227;
76: wave <=228;
77: wave <=229;
78: wave <=229;
79: wave <=230;
80: wave <=231;
81: wave <=232;
82: wave <=233;
83: wave <=234;
84: wave <=235;
85: wave <=235;
86: wave <=236;
87: wave <=237;
88: wave <=238;
89: wave <=239;
90: wave <=239;
91: wave <=240;
92: wave <=241;
93: wave <=241;
94: wave <=242;
95: wave <=243;
96: wave <=243;
97: wave <=244;
98: wave <=245;
99: wave <=245;
100: wave <=246;
101: wave <=246;
102: wave <=247;
103: wave <=247;
104: wave <=248;
105: wave <=248;
106: wave <=249;
107: wave <=249;
108: wave <=250;
109: wave <=250;
110: wave <=250;
111: wave <=251;
112: wave <=251;
113: wave <=251;
114: wave <=252;
115: wave <=252;
116: wave <=252;
117: wave <=253;
118: wave <=253;
119: wave <=253;
120: wave <=253;
121: wave <=254;
122: wave <=254;
123: wave <=254;
124: wave <=254;
125: wave <=254;
126: wave <=254;
127: wave <=254;
128: wave <=254;
129: wave <=254;
130: wave <=254;
131: wave <=254;
132: wave <=254;
133: wave <=254;
134: wave <=254;
135: wave <=254;
136: wave <=254;
137: wave <=254;
138: wave <=254;
139: wave <=254;
140: wave <=254;
141: wave <=254;
142: wave <=253;
143: wave <=253;
144: wave <=253;
145: wave <=253;
146: wave <=253;
147: wave <=252;
148: wave <=252;
149: wave <=252;
150: wave <=251;
151: wave <=251;
152: wave <=251;
153: wave <=250;
154: wave <=250;
155: wave <=249;
156: wave <=249;
157: wave <=248;
158: wave <=248;
159: wave <=248;
160: wave <=247;
161: wave <=247;
162: wave <=246;
163: wave <=245;
164: wave <=245;
165: wave <=244;
166: wave <=244;
167: wave <=243;
168: wave <=242;
169: wave <=242;
170: wave <=241;
171: wave <=240;
172: wave <=240;
173: wave <=239;
174: wave <=238;
175: wave <=237;
176: wave <=237;
177: wave <=236;
178: wave <=235;
179: wave <=234;
180: wave <=233;
181: wave <=233;
182: wave <=232;
183: wave <=231;
184: wave <=230;
185: wave <=229;
186: wave <=228;
187: wave <=227;
188: wave <=226;
189: wave <=225;
190: wave <=224;
191: wave <=223;
192: wave <=222;
193: wave <=221;
194: wave <=220;
195: wave <=219;
196: wave <=218;
197: wave <=217;
198: wave <=216;
199: wave <=215;
200: wave <=214;
201: wave <=213;
202: wave <=211;
203: wave <=210;
204: wave <=209;
205: wave <=208;
206: wave <=207;
207: wave <=206;
208: wave <=204;
209: wave <=203;
210: wave <=202;
211: wave <=201;
212: wave <=199;
213: wave <=198;
214: wave <=197;
215: wave <=196;
216: wave <=194;
217: wave <=193;
218: wave <=192;
219: wave <=190;
220: wave <=189;
221: wave <=188;
222: wave <=186;
223: wave <=185;
224: wave <=184;
225: wave <=182;
226: wave <=181;
227: wave <=180;
228: wave <=178;
229: wave <=177;
230: wave <=175;
231: wave <=174;
232: wave <=173;
233: wave <=171;
234: wave <=170;
235: wave <=168;
236: wave <=167;
237: wave <=165;
238: wave <=164;
239: wave <=162;
240: wave <=161;
241: wave <=159;
242: wave <=158;
243: wave <=156;
244: wave <=155;
245: wave <=154;
246: wave <=152;
247: wave <=151;
248: wave <=149;
249: wave <=148;
250: wave <=146;
251: wave <=144;
252: wave <=143;
253: wave <=141;
254: wave <=140;
255: wave <=138;
256: wave <=137;
257: wave <=135;
258: wave <=134;
259: wave <=132;
260: wave <=131;
261: wave <=129;
262: wave <=128;
263: wave <=126;
264: wave <=125;
265: wave <=123;
266: wave <=122;
267: wave <=120;
268: wave <=119;
269: wave <=117;
270: wave <=116;
271: wave <=114;
272: wave <=113;
273: wave <=111;
274: wave <=110;
275: wave <=108;
276: wave <=106;
277: wave <=105;
278: wave <=103;
279: wave <=102;
280: wave <=100;
281: wave <= 99;
282: wave <= 98;
283: wave <= 96;
284: wave <= 95;
285: wave <= 93;
286: wave <= 92;
287: wave <= 90;
288: wave <= 89;
289: wave <= 87;
290: wave <= 86;
291: wave <= 84;
292: wave <= 83;
293: wave <= 81;
294: wave <= 80;
295: wave <= 79;
296: wave <= 77;
297: wave <= 76;
298: wave <= 74;
299: wave <= 73;
300: wave <= 72;
301: wave <= 70;
302: wave <= 69;
303: wave <= 68;
304: wave <= 66;
305: wave <= 65;
306: wave <= 64;
307: wave <= 62;
308: wave <= 61;
309: wave <= 60;
310: wave <= 58;
311: wave <= 57;
312: wave <= 56;
313: wave <= 55;
314: wave <= 53;
315: wave <= 52;
316: wave <= 51;
317: wave <= 50;
318: wave <= 48;
319: wave <= 47;
320: wave <= 46;
321: wave <= 45;
322: wave <= 44;
323: wave <= 43;
324: wave <= 41;
325: wave <= 40;
326: wave <= 39;
327: wave <= 38;
328: wave <= 37;
329: wave <= 36;
330: wave <= 35;
331: wave <= 34;
332: wave <= 33;
333: wave <= 32;
334: wave <= 31;
335: wave <= 30;
336: wave <= 29;
337: wave <= 28;
338: wave <= 27;
339: wave <= 26;
340: wave <= 25;
341: wave <= 24;
342: wave <= 23;
343: wave <= 22;
344: wave <= 21;
345: wave <= 21;
346: wave <= 20;
347: wave <= 19;
348: wave <= 18;
349: wave <= 17;
350: wave <= 17;
351: wave <= 16;
352: wave <= 15;
353: wave <= 14;
354: wave <= 14;
355: wave <= 13;
356: wave <= 12;
357: wave <= 12;
358: wave <= 11;
359: wave <= 10;
360: wave <= 10;
361: wave <=  9;
362: wave <=  9;
363: wave <=  8;
364: wave <=  7;
365: wave <=  7;
366: wave <=  6;
367: wave <=  6;
368: wave <=  6;
369: wave <=  5;
370: wave <=  5;
371: wave <=  4;
372: wave <=  4;
373: wave <=  3;
374: wave <=  3;
375: wave <=  3;
376: wave <=  2;
377: wave <=  2;
378: wave <=  2;
379: wave <=  1;
380: wave <=  1;
381: wave <=  1;
382: wave <=  1;
383: wave <=  1;
384: wave <=  0;
385: wave <=  0;
386: wave <=  0;
387: wave <= -0;
388: wave <= -0;
389: wave <= -0;
390: wave <= -0;
391: wave <= -0;
392: wave <= -0;
393: wave <= -0;
394: wave <= -0;
395: wave <= -0;
396: wave <= -0;
397: wave <= -0;
398: wave <= -0;
399: wave <= -0;
400: wave <= -0;
401: wave <= -0;
402: wave <=  0;
403: wave <=  0;
404: wave <=  0;
405: wave <=  1;
406: wave <=  1;
407: wave <=  1;
408: wave <=  1;
409: wave <=  2;
410: wave <=  2;
411: wave <=  2;
412: wave <=  3;
413: wave <=  3;
414: wave <=  3;
415: wave <=  4;
416: wave <=  4;
417: wave <=  4;
418: wave <=  5;
419: wave <=  5;
420: wave <=  6;
421: wave <=  6;
422: wave <=  7;
423: wave <=  7;
424: wave <=  8;
425: wave <=  8;
426: wave <=  9;
427: wave <=  9;
428: wave <= 10;
429: wave <= 11;
430: wave <= 11;
431: wave <= 12;
432: wave <= 13;
433: wave <= 13;
434: wave <= 14;
435: wave <= 15;
436: wave <= 15;
437: wave <= 16;
438: wave <= 17;
439: wave <= 18;
440: wave <= 19;
441: wave <= 19;
442: wave <= 20;
443: wave <= 21;
444: wave <= 22;
445: wave <= 23;
446: wave <= 24;
447: wave <= 25;
448: wave <= 25;
449: wave <= 26;
450: wave <= 27;
451: wave <= 28;
452: wave <= 29;
453: wave <= 30;
454: wave <= 31;
455: wave <= 32;
456: wave <= 33;
457: wave <= 34;
458: wave <= 35;
459: wave <= 36;
460: wave <= 38;
461: wave <= 39;
462: wave <= 40;
463: wave <= 41;
464: wave <= 42;
465: wave <= 43;
466: wave <= 44;
467: wave <= 45;
468: wave <= 47;
469: wave <= 48;
470: wave <= 49;
471: wave <= 50;
472: wave <= 51;
473: wave <= 53;
474: wave <= 54;
475: wave <= 55;
476: wave <= 56;
477: wave <= 58;
478: wave <= 59;
479: wave <= 60;
480: wave <= 62;
481: wave <= 63;
482: wave <= 64;
483: wave <= 66;
484: wave <= 67;
485: wave <= 68;
486: wave <= 70;
487: wave <= 71;
488: wave <= 72;
489: wave <= 74;
490: wave <= 75;
491: wave <= 77;
492: wave <= 78;
493: wave <= 79;
494: wave <= 81;
495: wave <= 82;
496: wave <= 84;
497: wave <= 85;
498: wave <= 87;
499: wave <= 88;
500: wave <= 89;
501: wave <= 91;
502: wave <= 92;
503: wave <= 94;
504: wave <= 95;
505: wave <= 97;
506: wave <= 98;
507: wave <=100;
508: wave <=101;
509: wave <=103;
510: wave <=104;
511: wave <=106;
512: wave <=107;
513: wave <=109;
514: wave <=110;
515: wave <=112;
516: wave <=113;
517: wave <=115;
518: wave <=116;
519: wave <=118;
520: wave <=119;
521: wave <=121;
522: wave <=122;
523: wave <=124;
524: wave <=125;
	default: wave <= 127;
	endcase
end
endmodule
